`timescale 1ns / 1ps

module stat_machine(
    
);

endmodule