`timescale 1ns / 1ps

module calculate (
    input wire clk,
    input wire rst,
    input wire key_en,
    input wire equal,
    input wire [3: 0] in,
    output reg [15: 0] out
);

    


endmodule