`timescale 1ns / 1ps

module led ( 

);

endmodule