`timescale 1ns / 1ps

module keyboard( 
    
);

endmodule