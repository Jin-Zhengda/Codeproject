`timescale 1ns / 1ps

module state_machine(
    input wire clk,
    input wire rst,
    input wire en,
    input wire [3: 0] in,
    output reg [15: 0] result 
);




endmodule